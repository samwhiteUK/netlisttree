entity sub4 is
port map ();
subsub4b : entity work.another_submodule
port map ();

