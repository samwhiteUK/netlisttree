entity test_top_module is
sub1 : entity work.module
port map ();
sub2 : entity work.module
port map ();
sub3 : entity work.module
port map ();
sub4 : entity work.module
port map ();
sub5 : entity work.module
port map ();
sub6 : entity work.module
port map ();
sub7 : entity work.module
port map ();
sub8 : entity work.module
port map ();
sub9 : entity work.module2
port map ();
sub10 : entity work.module
port map ();
